module read_fifo(
    parameter integer ADDR_WIDTH = 64,
    parameter integer ID_WIDTH = 4,
    parameter integer DEPTH = 8
)(
    input logic clk,
    input logic rst_n,


);




endmodule